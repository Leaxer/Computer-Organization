module and_32bit (output [31:0] Y, input [31:0] A, input [31:0] B);
	and and1(Y[0], A[0], B[0]);
	and and2(Y[1], A[1], B[1]);
	and and3(Y[2], A[2], B[2]);
	and and4(Y[3], A[3], B[3]);
	and and5(Y[4], A[4], B[4]);
	and and6(Y[5], A[5], B[5]);
	and and7(Y[6], A[6], B[6]);
	and and8(Y[7], A[7], B[7]);
	and and9(Y[8], A[8], B[8]);
	and and10(Y[9], A[9], B[9]);
	and and11(Y[10], A[10], B[10]);
	and and12(Y[11], A[11], B[11]);
	and and13(Y[12], A[12], B[12]);
	and and14(Y[13], A[13], B[13]);
	and and15(Y[14], A[14], B[14]);
	and and16(Y[15], A[15], B[15]);
	and and17(Y[16], A[16], B[16]);
	and and18(Y[17], A[17], B[17]);
	and and19(Y[18], A[18], B[18]);
	and and20(Y[19], A[19], B[19]);
	and and21(Y[20], A[20], B[20]);
	and and22(Y[21], A[21], B[21]);
	and and23(Y[22], A[22], B[22]);
	and and24(Y[23], A[23], B[23]);
	and and25(Y[24], A[24], B[24]);
	and and26(Y[25], A[25], B[25]);
	and and27(Y[26], A[26], B[26]);
	and and28(Y[27], A[27], B[27]);
	and and29(Y[28], A[28], B[28]);
	and and30(Y[29], A[29], B[29]);
	and and31(Y[30], A[30], B[30]);
	and and32(Y[31], A[31], B[31]);
endmodule
module xor_32bit (output [31:0] Y, input [31:0] A, input [31:0] B);
	xor xor1(Y[0], A[0], B[0]);
	xor xor2(Y[1], A[1], B[1]);
	xor xor3(Y[2], A[2], B[2]);
	xor xor4(Y[3], A[3], B[3]);
	xor xor5(Y[4], A[4], B[4]);
	xor xor6(Y[5], A[5], B[5]);
	xor xor7(Y[6], A[6], B[6]);
	xor xor8(Y[7], A[7], B[7]);
	xor xor9(Y[8], A[8], B[8]);
	xor xor10(Y[9], A[9] ,B[9]);
	xor xor11(Y[10], A[10], B[10]);
	xor xor12(Y[11], A[11], B[11]);
	xor xor13(Y[12], A[12], B[12]);
	xor xor14(Y[13], A[13], B[13]);
	xor xor15(Y[14], A[14], B[14]);
	xor xor16(Y[15], A[15], B[15]);
	xor xor17(Y[16], A[16], B[16]);
	xor xor18(Y[17], A[17], B[17]);
	xor xor19(Y[18], A[18], B[18]);
	xor xor20(Y[19], A[19], B[19]);
	xor xor21(Y[20], A[20], B[20]);
	xor xor22(Y[21], A[21], B[21]);
	xor xor23(Y[22], A[22], B[22]);
	xor xor24(Y[23], A[23], B[23]);
	xor xor25(Y[24], A[24], B[24]);
	xor xor26(Y[25], A[25], B[25]);
	xor xor27(Y[26], A[26], B[26]);
	xor xor28(Y[27], A[27], B[27]);
	xor xor29(Y[28], A[28], B[28]);
	xor xor30(Y[29], A[29], B[29]);
	xor xor31(Y[30], A[30], B[30]);
	xor xor32(Y[31], A[31], B[31]);
endmodule

module sign_extend (output [31:0] sign_ext_imm, input [15:0] imm);
   or or1(sign_ext_imm[0], 1'b0, imm[0]);
	or or2(sign_ext_imm[1], 1'b0, imm[1]);
	or or3(sign_ext_imm[2], 1'b0, imm[2]);
	or or4(sign_ext_imm[3], 1'b0, imm[3]);
	or or5(sign_ext_imm[4], 1'b0, imm[4]);
	or or6(sign_ext_imm[5], 1'b0, imm[5]);
	or or7(sign_ext_imm[6], 1'b0, imm[6]);
	or or8(sign_ext_imm[7], 1'b0, imm[7]);
	or or9(sign_ext_imm[8], 1'b0, imm[8]);
	or or10(sign_ext_imm[9], 1'b0, imm[9]);
	or or11(sign_ext_imm[10], 1'b0, imm[10]);
	or or12(sign_ext_imm[11], 1'b0, imm[11]);
	or or13(sign_ext_imm[12], 1'b0, imm[12]);
	or or14(sign_ext_imm[13], 1'b0, imm[13]);
	or or15(sign_ext_imm[14], 1'b0, imm[14]);
	or or16(sign_ext_imm[15], 1'b0, imm[15]);
	and and1(sign_ext_imm[16], 1'b1, imm[15]);
	and and2(sign_ext_imm[17], 1'b1, imm[15]);
	and and3(sign_ext_imm[18], 1'b1, imm[15]);
	and and4(sign_ext_imm[19], 1'b1, imm[15]);
	and and5(sign_ext_imm[20], 1'b1, imm[15]);
	and and6(sign_ext_imm[21], 1'b1, imm[15]);
	and and7(sign_ext_imm[22], 1'b1, imm[15]);
	and and8(sign_ext_imm[23], 1'b1, imm[15]);
	and and9(sign_ext_imm[24], 1'b1, imm[15]);
	and and10(sign_ext_imm[25], 1'b1, imm[15]);
	and and11(sign_ext_imm[26], 1'b1, imm[15]);
	and and12(sign_ext_imm[27], 1'b1, imm[15]);
	and and13(sign_ext_imm[28], 1'b1, imm[15]);
	and and14(sign_ext_imm[29], 1'b1, imm[15]);
	and and15(sign_ext_imm[30], 1'b1, imm[15]);
	and and16(sign_ext_imm[31], 1'b1, imm[15]);

endmodule
module sign_extend_alu32bit (output [31:0] Y, input x);
	and and1(Y[0], 1'b1, x);
	and and2(Y[1], 1'b1, x);
	and and3(Y[2], 1'b1, x);
	and and4(Y[3], 1'b1, x);
	and and5(Y[4], 1'b1, x);
	and and6(Y[5], 1'b1, x);
	and and7(Y[6], 1'b1, x);
	and and8(Y[7], 1'b1, x);
	and and9(Y[8], 1'b1, x);
	and and10(Y[9], 1'b1, x);
	and and11(Y[10], 1'b1, x);
	and and12(Y[11], 1'b1, x);
	and and13(Y[12], 1'b1, x);
	and and14(Y[13], 1'b1, x);
	and and15(Y[14], 1'b1, x);
	and and16(Y[15], 1'b1, x);
	and and17(Y[16], 1'b1, x);
	and and18(Y[17], 1'b1, x);
	and and19(Y[18], 1'b1, x);
	and and20(Y[19], 1'b1, x);
	and and21(Y[20], 1'b1, x);
	and and22(Y[21], 1'b1, x);
	and and23(Y[22], 1'b1, x);
	and and24(Y[23], 1'b1, x);
	and and25(Y[24], 1'b1, x);
	and and26(Y[25], 1'b1, x);
	and and27(Y[26], 1'b1, x);
	and and28(Y[27], 1'b1, x);
	and and29(Y[28], 1'b1, x);
	and and30(Y[29], 1'b1, x);
	and and31(Y[30], 1'b1, x);
	and and32(Y[31], 1'b1, x);
endmodule
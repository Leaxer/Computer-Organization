module buf_32bit (output [31:0] Y, input [31:0] X);
	buf buf1(Y[0], X[0]);
	buf buf2(Y[1], X[1]);
	buf buf3(Y[2], X[2]);
	buf buf4(Y[3], X[3]);
	buf buf5(Y[4], X[4]);
	buf buf6(Y[5], X[5]);
	buf buf7(Y[6], X[6]);
	buf buf8(Y[7], X[7]);
	buf buf9(Y[8], X[8]);
	buf buf10(Y[9], X[9]);
	buf buf11(Y[10], X[10]);
	buf buf12(Y[11], X[11]);
	buf buf13(Y[12], X[12]);
	buf buf14(Y[13], X[13]);
	buf buf15(Y[14], X[14]);
	buf buf16(Y[15], X[15]);
	buf buf17(Y[16], X[16]);
	buf buf18(Y[17], X[17]);
	buf buf19(Y[18], X[18]);
	buf buf20(Y[19], X[19]);
	buf buf21(Y[20], X[20]);
	buf buf22(Y[21], X[21]);
	buf buf23(Y[22], X[22]);
	buf buf24(Y[23], X[23]);
	buf buf25(Y[24], X[24]);
	buf buf26(Y[25], X[25]);
	buf buf27(Y[26], X[26]);
	buf buf28(Y[27], X[27]);
	buf buf29(Y[28], X[28]);
	buf buf30(Y[29], X[29]);
	buf buf31(Y[30], X[30]);
	buf buf32(Y[31], X[31]);
endmodule
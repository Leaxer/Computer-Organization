module nor_32bit (output [31:0] Y, input [31:0] A, input [31:0] B);
	nor nor1(Y[0], A[0], B[0]);
	nor nor2(Y[1], A[1], B[1]);
	nor nor3(Y[2], A[2], B[2]);
	nor nor4(Y[3], A[3], B[3]);
	nor nor5(Y[4], A[4], B[4]);
	nor nor6(Y[5], A[5], B[5]);
	nor nor7(Y[6], A[6], B[6]);
	nor nor8(Y[7], A[7], B[7]);
	nor nor9(Y[8], A[8], B[8]);
	nor nor10(Y[9], A[9] ,B[9]);
	nor nor11(Y[10], A[10], B[10]);
	nor nor12(Y[11], A[11], B[11]);
	nor nor13(Y[12], A[12], B[12]);
	nor nor14(Y[13], A[13], B[13]);
	nor nor15(Y[14], A[14], B[14]);
	nor nor16(Y[15], A[15], B[15]);
	nor nor17(Y[16], A[16], B[16]);
	nor nor18(Y[17], A[17], B[17]);
	nor nor19(Y[18], A[18], B[18]);
	nor nor20(Y[19], A[19], B[19]);
	nor nor21(Y[20], A[20], B[20]);
	nor nor22(Y[21], A[21], B[21]);
	nor nor23(Y[22], A[22], B[22]);
	nor nor24(Y[23], A[23], B[23]);
	nor nor25(Y[24], A[24], B[24]);
	nor nor26(Y[25], A[25], B[25]);
	nor nor27(Y[26], A[26], B[26]);
	nor nor28(Y[27], A[27], B[27]);
	nor nor29(Y[28], A[28], B[28]);
	nor nor30(Y[29], A[29], B[29]);
	nor nor31(Y[30], A[30], B[30]);
	nor nor32(Y[31], A[31], B[31]);
endmodule